parameter ALU_OP_WIDTH = 6,
parameter N_HWLP      = 1,
parameter N_HWLP_BITS = $clog2(N_HWLP),
parameter DBG_SETS_W = 6,
parameter RDATA_WIDTH = 32,
parameter N_EXT_CNT    = 0,
parameter N_EXT_PERF_COUNTERS = 0,
parameter INSTR_RDATA_WIDTH   = 32
