parameter ALU_OP_WIDTH = 6,
parameter DBG_SETS_W = 6
