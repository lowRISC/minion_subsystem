parameter ALU_OP_WIDTH = 6,
parameter DBG_SETS_W = 6,
parameter RDATA_WIDTH = 32,
parameter N_EXT_CNT    = 0,
parameter N_EXT_PERF_COUNTERS = 0,
parameter INSTR_RDATA_WIDTH   = 32
