module clk_wiz_arty_0
 (
 // Clock in ports
  input         clk_in1,
  // Clock out ports
  output        msoc_clk
 );

 assign msoc_clk = clk_in1;

endmodule

module ila_arty_0 (
clk,


probe0,
probe1,
probe2,
probe3,
probe4,
probe5,
probe6,
probe7,
probe8,
probe9,
probe10,
probe11,
probe12,
probe13
);

input clk;


input [0 : 0] probe0;
input [0 : 0] probe1;
input [0 : 0] probe2;
input [31 : 0] probe3;
input [31 : 0] probe4;
input [0 : 0] probe5;
input [3 : 0] probe6;
input [0 : 0] probe7;
input [7 : 0] probe8;
input [0 : 0] probe9;
input [15 : 0] probe10;
input [31 : 0] probe11;
input [0 : 0] probe12;
input [3 : 0] probe13;

endmodule
