module dpram(clka, clkb, dina, addra, wea, douta, ena, dinb, addrb, web, doutb, enb);

   parameter rwidth = 14;

   input clka;
   input clkb;
   input [127:0] dina;
   input [13:0]  addra;
   input [0:0]   wea;
   input [15:0]  ena;
   output [127:0] douta;
   input [127:0]  dinb;
   input [13:0]   addrb;
   input [0:0]    web;
   input [15:0]   enb;
   output [127:0] doutb;

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_0 (
                                               .CLKA(clka),      // Port A Clock
                                               .DOA(douta[0]),  // Port A 1-bit Data Output
                                               .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                               .DIA(dina[0]),   // Port A 1-bit Data Input
                                               .ENA(ena[0]),    // Port A RAM Enable Input
                                               .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                               .WEA(wea),         // Port A Write Enable Input
                                               .CLKB(clkb),      // Port B Clock
                                               .DOB(doutb[0]),  // Port B 1-bit Data Output
                                               .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                               .DIB(dinb[0]),   // Port B 1-bit Data Input
                                               .ENB(enb[0]),    // Port B RAM Enable Input
                                               .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                               .WEB(web)         // Port B Write Enable Input
                                               ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_1 (
                                               .CLKA(clka),      // Port A Clock
                                               .DOA(douta[1]),  // Port A 1-bit Data Output
                                               .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                               .DIA(dina[1]),   // Port A 1-bit Data Input
                                               .ENA(ena[0]),    // Port A RAM Enable Input
                                               .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                               .WEA(wea),         // Port A Write Enable Input
                                               .CLKB(clkb),      // Port B Clock
                                               .DOB(doutb[1]),  // Port B 1-bit Data Output
                                               .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                               .DIB(dinb[1]),   // Port B 1-bit Data Input
                                               .ENB(enb[0]),    // Port B RAM Enable Input
                                               .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                               .WEB(web)         // Port B Write Enable Input
                                               ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_2 (
                                               .CLKA(clka),      // Port A Clock
                                               .DOA(douta[2]),  // Port A 1-bit Data Output
                                               .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                               .DIA(dina[2]),   // Port A 1-bit Data Input
                                               .ENA(ena[0]),    // Port A RAM Enable Input
                                               .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                               .WEA(wea),         // Port A Write Enable Input
                                               .CLKB(clkb),      // Port B Clock
                                               .DOB(doutb[2]),  // Port B 1-bit Data Output
                                               .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                               .DIB(dinb[2]),   // Port B 1-bit Data Input
                                               .ENB(enb[0]),    // Port B RAM Enable Input
                                               .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                               .WEB(web)         // Port B Write Enable Input
                                               ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_3 (
                                               .CLKA(clka),      // Port A Clock
                                               .DOA(douta[3]),  // Port A 1-bit Data Output
                                               .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                               .DIA(dina[3]),   // Port A 1-bit Data Input
                                               .ENA(ena[0]),    // Port A RAM Enable Input
                                               .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                               .WEA(wea),         // Port A Write Enable Input
                                               .CLKB(clkb),      // Port B Clock
                                               .DOB(doutb[3]),  // Port B 1-bit Data Output
                                               .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                               .DIB(dinb[3]),   // Port B 1-bit Data Input
                                               .ENB(enb[0]),    // Port B RAM Enable Input
                                               .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                               .WEB(web)         // Port B Write Enable Input
                                               ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_4 (
                                               .CLKA(clka),      // Port A Clock
                                               .DOA(douta[4]),  // Port A 1-bit Data Output
                                               .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                               .DIA(dina[4]),   // Port A 1-bit Data Input
                                               .ENA(ena[0]),    // Port A RAM Enable Input
                                               .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                               .WEA(wea),         // Port A Write Enable Input
                                               .CLKB(clkb),      // Port B Clock
                                               .DOB(doutb[4]),  // Port B 1-bit Data Output
                                               .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                               .DIB(dinb[4]),   // Port B 1-bit Data Input
                                               .ENB(enb[0]),    // Port B RAM Enable Input
                                               .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                               .WEB(web)         // Port B Write Enable Input
                                               ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_5 (
                                               .CLKA(clka),      // Port A Clock
                                               .DOA(douta[5]),  // Port A 1-bit Data Output
                                               .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                               .DIA(dina[5]),   // Port A 1-bit Data Input
                                               .ENA(ena[0]),    // Port A RAM Enable Input
                                               .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                               .WEA(wea),         // Port A Write Enable Input
                                               .CLKB(clkb),      // Port B Clock
                                               .DOB(doutb[5]),  // Port B 1-bit Data Output
                                               .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                               .DIB(dinb[5]),   // Port B 1-bit Data Input
                                               .ENB(enb[0]),    // Port B RAM Enable Input
                                               .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                               .WEB(web)         // Port B Write Enable Input
                                               ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_6 (
                                               .CLKA(clka),      // Port A Clock
                                               .DOA(douta[6]),  // Port A 1-bit Data Output
                                               .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                               .DIA(dina[6]),   // Port A 1-bit Data Input
                                               .ENA(ena[0]),    // Port A RAM Enable Input
                                               .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                               .WEA(wea),         // Port A Write Enable Input
                                               .CLKB(clkb),      // Port B Clock
                                               .DOB(doutb[6]),  // Port B 1-bit Data Output
                                               .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                               .DIB(dinb[6]),   // Port B 1-bit Data Input
                                               .ENB(enb[0]),    // Port B RAM Enable Input
                                               .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                               .WEB(web)         // Port B Write Enable Input
                                               ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_7 (
                                               .CLKA(clka),      // Port A Clock
                                               .DOA(douta[7]),  // Port A 1-bit Data Output
                                               .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                               .DIA(dina[7]),   // Port A 1-bit Data Input
                                               .ENA(ena[0]),    // Port A RAM Enable Input
                                               .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                               .WEA(wea),         // Port A Write Enable Input
                                               .CLKB(clkb),      // Port B Clock
                                               .DOB(doutb[7]),  // Port B 1-bit Data Output
                                               .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                               .DIB(dinb[7]),   // Port B 1-bit Data Input
                                               .ENB(enb[0]),    // Port B RAM Enable Input
                                               .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                               .WEB(web)         // Port B Write Enable Input
                                               ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_8 (
                                               .CLKA(clka),      // Port A Clock
                                               .DOA(douta[8]),  // Port A 1-bit Data Output
                                               .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                               .DIA(dina[8]),   // Port A 1-bit Data Input
                                               .ENA(ena[1]),    // Port A RAM Enable Input
                                               .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                               .WEA(wea),         // Port A Write Enable Input
                                               .CLKB(clkb),      // Port B Clock
                                               .DOB(doutb[8]),  // Port B 1-bit Data Output
                                               .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                               .DIB(dinb[8]),   // Port B 1-bit Data Input
                                               .ENB(enb[1]),    // Port B RAM Enable Input
                                               .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                               .WEB(web)         // Port B Write Enable Input
                                               ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_9 (
                                               .CLKA(clka),      // Port A Clock
                                               .DOA(douta[9]),  // Port A 1-bit Data Output
                                               .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                               .DIA(dina[9]),   // Port A 1-bit Data Input
                                               .ENA(ena[1]),    // Port A RAM Enable Input
                                               .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                               .WEA(wea),         // Port A Write Enable Input
                                               .CLKB(clkb),      // Port B Clock
                                               .DOB(doutb[9]),  // Port B 1-bit Data Output
                                               .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                               .DIB(dinb[9]),   // Port B 1-bit Data Input
                                               .ENB(enb[1]),    // Port B RAM Enable Input
                                               .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                               .WEB(web)         // Port B Write Enable Input
                                               ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_10 (
                                                .CLKA(clka),      // Port A Clock
                                                .DOA(douta[10]),  // Port A 1-bit Data Output
                                                .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                .DIA(dina[10]),   // Port A 1-bit Data Input
                                                .ENA(ena[1]),    // Port A RAM Enable Input
                                                .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                .WEA(wea),         // Port A Write Enable Input
                                                .CLKB(clkb),      // Port B Clock
                                                .DOB(doutb[10]),  // Port B 1-bit Data Output
                                                .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                .DIB(dinb[10]),   // Port B 1-bit Data Input
                                                .ENB(enb[1]),    // Port B RAM Enable Input
                                                .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                .WEB(web)         // Port B Write Enable Input
                                                ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_11 (
                                                .CLKA(clka),      // Port A Clock
                                                .DOA(douta[11]),  // Port A 1-bit Data Output
                                                .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                .DIA(dina[11]),   // Port A 1-bit Data Input
                                                .ENA(ena[1]),    // Port A RAM Enable Input
                                                .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                .WEA(wea),         // Port A Write Enable Input
                                                .CLKB(clkb),      // Port B Clock
                                                .DOB(doutb[11]),  // Port B 1-bit Data Output
                                                .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                .DIB(dinb[11]),   // Port B 1-bit Data Input
                                                .ENB(enb[1]),    // Port B RAM Enable Input
                                                .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                .WEB(web)         // Port B Write Enable Input
                                                ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_12 (
                                                .CLKA(clka),      // Port A Clock
                                                .DOA(douta[12]),  // Port A 1-bit Data Output
                                                .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                .DIA(dina[12]),   // Port A 1-bit Data Input
                                                .ENA(ena[1]),    // Port A RAM Enable Input
                                                .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                .WEA(wea),         // Port A Write Enable Input
                                                .CLKB(clkb),      // Port B Clock
                                                .DOB(doutb[12]),  // Port B 1-bit Data Output
                                                .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                .DIB(dinb[12]),   // Port B 1-bit Data Input
                                                .ENB(enb[1]),    // Port B RAM Enable Input
                                                .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                .WEB(web)         // Port B Write Enable Input
                                                ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_13 (
                                                .CLKA(clka),      // Port A Clock
                                                .DOA(douta[13]),  // Port A 1-bit Data Output
                                                .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                .DIA(dina[13]),   // Port A 1-bit Data Input
                                                .ENA(ena[1]),    // Port A RAM Enable Input
                                                .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                .WEA(wea),         // Port A Write Enable Input
                                                .CLKB(clkb),      // Port B Clock
                                                .DOB(doutb[13]),  // Port B 1-bit Data Output
                                                .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                .DIB(dinb[13]),   // Port B 1-bit Data Input
                                                .ENB(enb[1]),    // Port B RAM Enable Input
                                                .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                .WEB(web)         // Port B Write Enable Input
                                                ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_14 (
                                                .CLKA(clka),      // Port A Clock
                                                .DOA(douta[14]),  // Port A 1-bit Data Output
                                                .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                .DIA(dina[14]),   // Port A 1-bit Data Input
                                                .ENA(ena[1]),    // Port A RAM Enable Input
                                                .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                .WEA(wea),         // Port A Write Enable Input
                                                .CLKB(clkb),      // Port B Clock
                                                .DOB(doutb[14]),  // Port B 1-bit Data Output
                                                .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                .DIB(dinb[14]),   // Port B 1-bit Data Input
                                                .ENB(enb[1]),    // Port B RAM Enable Input
                                                .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                .WEB(web)         // Port B Write Enable Input
                                                ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_15 (
                                                .CLKA(clka),      // Port A Clock
                                                .DOA(douta[15]),  // Port A 1-bit Data Output
                                                .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                .DIA(dina[15]),   // Port A 1-bit Data Input
                                                .ENA(ena[1]),    // Port A RAM Enable Input
                                                .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                .WEA(wea),         // Port A Write Enable Input
                                                .CLKB(clkb),      // Port B Clock
                                                .DOB(doutb[15]),  // Port B 1-bit Data Output
                                                .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                .DIB(dinb[15]),   // Port B 1-bit Data Input
                                                .ENB(enb[1]),    // Port B RAM Enable Input
                                                .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                .WEB(web)         // Port B Write Enable Input
                                                ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_16 (
                                                .CLKA(clka),      // Port A Clock
                                                .DOA(douta[16]),  // Port A 1-bit Data Output
                                                .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                .DIA(dina[16]),   // Port A 1-bit Data Input
                                                .ENA(ena[2]),    // Port A RAM Enable Input
                                                .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                .WEA(wea),         // Port A Write Enable Input
                                                .CLKB(clkb),      // Port B Clock
                                                .DOB(doutb[16]),  // Port B 1-bit Data Output
                                                .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                .DIB(dinb[16]),   // Port B 1-bit Data Input
                                                .ENB(enb[2]),    // Port B RAM Enable Input
                                                .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                .WEB(web)         // Port B Write Enable Input
                                                ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_17 (
                                                .CLKA(clka),      // Port A Clock
                                                .DOA(douta[17]),  // Port A 1-bit Data Output
                                                .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                .DIA(dina[17]),   // Port A 1-bit Data Input
                                                .ENA(ena[2]),    // Port A RAM Enable Input
                                                .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                .WEA(wea),         // Port A Write Enable Input
                                                .CLKB(clkb),      // Port B Clock
                                                .DOB(doutb[17]),  // Port B 1-bit Data Output
                                                .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                .DIB(dinb[17]),   // Port B 1-bit Data Input
                                                .ENB(enb[2]),    // Port B RAM Enable Input
                                                .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                .WEB(web)         // Port B Write Enable Input
                                                ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_18 (
                                                .CLKA(clka),      // Port A Clock
                                                .DOA(douta[18]),  // Port A 1-bit Data Output
                                                .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                .DIA(dina[18]),   // Port A 1-bit Data Input
                                                .ENA(ena[2]),    // Port A RAM Enable Input
                                                .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                .WEA(wea),         // Port A Write Enable Input
                                                .CLKB(clkb),      // Port B Clock
                                                .DOB(doutb[18]),  // Port B 1-bit Data Output
                                                .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                .DIB(dinb[18]),   // Port B 1-bit Data Input
                                                .ENB(enb[2]),    // Port B RAM Enable Input
                                                .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                .WEB(web)         // Port B Write Enable Input
                                                ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_19 (
                                                .CLKA(clka),      // Port A Clock
                                                .DOA(douta[19]),  // Port A 1-bit Data Output
                                                .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                .DIA(dina[19]),   // Port A 1-bit Data Input
                                                .ENA(ena[2]),    // Port A RAM Enable Input
                                                .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                .WEA(wea),         // Port A Write Enable Input
                                                .CLKB(clkb),      // Port B Clock
                                                .DOB(doutb[19]),  // Port B 1-bit Data Output
                                                .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                .DIB(dinb[19]),   // Port B 1-bit Data Input
                                                .ENB(enb[2]),    // Port B RAM Enable Input
                                                .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                .WEB(web)         // Port B Write Enable Input
                                                ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_20 (
                                                .CLKA(clka),      // Port A Clock
                                                .DOA(douta[20]),  // Port A 1-bit Data Output
                                                .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                .DIA(dina[20]),   // Port A 1-bit Data Input
                                                .ENA(ena[2]),    // Port A RAM Enable Input
                                                .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                .WEA(wea),         // Port A Write Enable Input
                                                .CLKB(clkb),      // Port B Clock
                                                .DOB(doutb[20]),  // Port B 1-bit Data Output
                                                .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                .DIB(dinb[20]),   // Port B 1-bit Data Input
                                                .ENB(enb[2]),    // Port B RAM Enable Input
                                                .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                .WEB(web)         // Port B Write Enable Input
                                                ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_21 (
                                                .CLKA(clka),      // Port A Clock
                                                .DOA(douta[21]),  // Port A 1-bit Data Output
                                                .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                .DIA(dina[21]),   // Port A 1-bit Data Input
                                                .ENA(ena[2]),    // Port A RAM Enable Input
                                                .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                .WEA(wea),         // Port A Write Enable Input
                                                .CLKB(clkb),      // Port B Clock
                                                .DOB(doutb[21]),  // Port B 1-bit Data Output
                                                .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                .DIB(dinb[21]),   // Port B 1-bit Data Input
                                                .ENB(enb[2]),    // Port B RAM Enable Input
                                                .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                .WEB(web)         // Port B Write Enable Input
                                                ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_22 (
                                                .CLKA(clka),      // Port A Clock
                                                .DOA(douta[22]),  // Port A 1-bit Data Output
                                                .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                .DIA(dina[22]),   // Port A 1-bit Data Input
                                                .ENA(ena[2]),    // Port A RAM Enable Input
                                                .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                .WEA(wea),         // Port A Write Enable Input
                                                .CLKB(clkb),      // Port B Clock
                                                .DOB(doutb[22]),  // Port B 1-bit Data Output
                                                .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                .DIB(dinb[22]),   // Port B 1-bit Data Input
                                                .ENB(enb[2]),    // Port B RAM Enable Input
                                                .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                .WEB(web)         // Port B Write Enable Input
                                                ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_23 (
                                                .CLKA(clka),      // Port A Clock
                                                .DOA(douta[23]),  // Port A 1-bit Data Output
                                                .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                .DIA(dina[23]),   // Port A 1-bit Data Input
                                                .ENA(ena[2]),    // Port A RAM Enable Input
                                                .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                .WEA(wea),         // Port A Write Enable Input
                                                .CLKB(clkb),      // Port B Clock
                                                .DOB(doutb[23]),  // Port B 1-bit Data Output
                                                .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                .DIB(dinb[23]),   // Port B 1-bit Data Input
                                                .ENB(enb[2]),    // Port B RAM Enable Input
                                                .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                .WEB(web)         // Port B Write Enable Input
                                                ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_24 (
                                                .CLKA(clka),      // Port A Clock
                                                .DOA(douta[24]),  // Port A 1-bit Data Output
                                                .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                .DIA(dina[24]),   // Port A 1-bit Data Input
                                                .ENA(ena[3]),    // Port A RAM Enable Input
                                                .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                .WEA(wea),         // Port A Write Enable Input
                                                .CLKB(clkb),      // Port B Clock
                                                .DOB(doutb[24]),  // Port B 1-bit Data Output
                                                .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                .DIB(dinb[24]),   // Port B 1-bit Data Input
                                                .ENB(enb[3]),    // Port B RAM Enable Input
                                                .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                .WEB(web)         // Port B Write Enable Input
                                                ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_25 (
                                                .CLKA(clka),      // Port A Clock
                                                .DOA(douta[25]),  // Port A 1-bit Data Output
                                                .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                .DIA(dina[25]),   // Port A 1-bit Data Input
                                                .ENA(ena[3]),    // Port A RAM Enable Input
                                                .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                .WEA(wea),         // Port A Write Enable Input
                                                .CLKB(clkb),      // Port B Clock
                                                .DOB(doutb[25]),  // Port B 1-bit Data Output
                                                .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                .DIB(dinb[25]),   // Port B 1-bit Data Input
                                                .ENB(enb[3]),    // Port B RAM Enable Input
                                                .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                .WEB(web)         // Port B Write Enable Input
                                                ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_26 (
                                                .CLKA(clka),      // Port A Clock
                                                .DOA(douta[26]),  // Port A 1-bit Data Output
                                                .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                .DIA(dina[26]),   // Port A 1-bit Data Input
                                                .ENA(ena[3]),    // Port A RAM Enable Input
                                                .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                .WEA(wea),         // Port A Write Enable Input
                                                .CLKB(clkb),      // Port B Clock
                                                .DOB(doutb[26]),  // Port B 1-bit Data Output
                                                .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                .DIB(dinb[26]),   // Port B 1-bit Data Input
                                                .ENB(enb[3]),    // Port B RAM Enable Input
                                                .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                .WEB(web)         // Port B Write Enable Input
                                                ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_27 (
                                                .CLKA(clka),      // Port A Clock
                                                .DOA(douta[27]),  // Port A 1-bit Data Output
                                                .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                .DIA(dina[27]),   // Port A 1-bit Data Input
                                                .ENA(ena[3]),    // Port A RAM Enable Input
                                                .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                .WEA(wea),         // Port A Write Enable Input
                                                .CLKB(clkb),      // Port B Clock
                                                .DOB(doutb[27]),  // Port B 1-bit Data Output
                                                .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                .DIB(dinb[27]),   // Port B 1-bit Data Input
                                                .ENB(enb[3]),    // Port B RAM Enable Input
                                                .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                .WEB(web)         // Port B Write Enable Input
                                                ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_28 (
                                                .CLKA(clka),      // Port A Clock
                                                .DOA(douta[28]),  // Port A 1-bit Data Output
                                                .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                .DIA(dina[28]),   // Port A 1-bit Data Input
                                                .ENA(ena[3]),    // Port A RAM Enable Input
                                                .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                .WEA(wea),         // Port A Write Enable Input
                                                .CLKB(clkb),      // Port B Clock
                                                .DOB(doutb[28]),  // Port B 1-bit Data Output
                                                .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                .DIB(dinb[28]),   // Port B 1-bit Data Input
                                                .ENB(enb[3]),    // Port B RAM Enable Input
                                                .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                .WEB(web)         // Port B Write Enable Input
                                                ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_29 (
                                                .CLKA(clka),      // Port A Clock
                                                .DOA(douta[29]),  // Port A 1-bit Data Output
                                                .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                .DIA(dina[29]),   // Port A 1-bit Data Input
                                                .ENA(ena[3]),    // Port A RAM Enable Input
                                                .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                .WEA(wea),         // Port A Write Enable Input
                                                .CLKB(clkb),      // Port B Clock
                                                .DOB(doutb[29]),  // Port B 1-bit Data Output
                                                .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                .DIB(dinb[29]),   // Port B 1-bit Data Input
                                                .ENB(enb[3]),    // Port B RAM Enable Input
                                                .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                .WEB(web)         // Port B Write Enable Input
                                                ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_30 (
                                                .CLKA(clka),      // Port A Clock
                                                .DOA(douta[30]),  // Port A 1-bit Data Output
                                                .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                .DIA(dina[30]),   // Port A 1-bit Data Input
                                                .ENA(ena[3]),    // Port A RAM Enable Input
                                                .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                .WEA(wea),         // Port A Write Enable Input
                                                .CLKB(clkb),      // Port B Clock
                                                .DOB(doutb[30]),  // Port B 1-bit Data Output
                                                .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                .DIB(dinb[30]),   // Port B 1-bit Data Input
                                                .ENB(enb[3]),    // Port B RAM Enable Input
                                                .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                .WEB(web)         // Port B Write Enable Input
                                                ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_31 (
                                                .CLKA(clka),      // Port A Clock
                                                .DOA(douta[31]),  // Port A 1-bit Data Output
                                                .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                .DIA(dina[31]),   // Port A 1-bit Data Input
                                                .ENA(ena[3]),    // Port A RAM Enable Input
                                                .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                .WEA(wea),         // Port A Write Enable Input
                                                .CLKB(clkb),      // Port B Clock
                                                .DOB(doutb[31]),  // Port B 1-bit Data Output
                                                .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                .DIB(dinb[31]),   // Port B 1-bit Data Input
                                                .ENB(enb[3]),    // Port B RAM Enable Input
                                                .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                .WEB(web)         // Port B Write Enable Input
                                                ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_32 (
                                                .CLKA(clka),      // Port A Clock
                                                .DOA(douta[32]),  // Port A 1-bit Data Output
                                                .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                .DIA(dina[32]),   // Port A 1-bit Data Input
                                                .ENA(ena[4]),    // Port A RAM Enable Input
                                                .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                .WEA(wea),         // Port A Write Enable Input
                                                .CLKB(clkb),      // Port B Clock
                                                .DOB(doutb[32]),  // Port B 1-bit Data Output
                                                .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                .DIB(dinb[32]),   // Port B 1-bit Data Input
                                                .ENB(enb[4]),    // Port B RAM Enable Input
                                                .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                .WEB(web)         // Port B Write Enable Input
                                                ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_33 (
                                                .CLKA(clka),      // Port A Clock
                                                .DOA(douta[33]),  // Port A 1-bit Data Output
                                                .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                .DIA(dina[33]),   // Port A 1-bit Data Input
                                                .ENA(ena[4]),    // Port A RAM Enable Input
                                                .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                .WEA(wea),         // Port A Write Enable Input
                                                .CLKB(clkb),      // Port B Clock
                                                .DOB(doutb[33]),  // Port B 1-bit Data Output
                                                .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                .DIB(dinb[33]),   // Port B 1-bit Data Input
                                                .ENB(enb[4]),    // Port B RAM Enable Input
                                                .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                .WEB(web)         // Port B Write Enable Input
                                                ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_34 (
                                                .CLKA(clka),      // Port A Clock
                                                .DOA(douta[34]),  // Port A 1-bit Data Output
                                                .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                .DIA(dina[34]),   // Port A 1-bit Data Input
                                                .ENA(ena[4]),    // Port A RAM Enable Input
                                                .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                .WEA(wea),         // Port A Write Enable Input
                                                .CLKB(clkb),      // Port B Clock
                                                .DOB(doutb[34]),  // Port B 1-bit Data Output
                                                .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                .DIB(dinb[34]),   // Port B 1-bit Data Input
                                                .ENB(enb[4]),    // Port B RAM Enable Input
                                                .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                .WEB(web)         // Port B Write Enable Input
                                                ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_35 (
                                                .CLKA(clka),      // Port A Clock
                                                .DOA(douta[35]),  // Port A 1-bit Data Output
                                                .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                .DIA(dina[35]),   // Port A 1-bit Data Input
                                                .ENA(ena[4]),    // Port A RAM Enable Input
                                                .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                .WEA(wea),         // Port A Write Enable Input
                                                .CLKB(clkb),      // Port B Clock
                                                .DOB(doutb[35]),  // Port B 1-bit Data Output
                                                .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                .DIB(dinb[35]),   // Port B 1-bit Data Input
                                                .ENB(enb[4]),    // Port B RAM Enable Input
                                                .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                .WEB(web)         // Port B Write Enable Input
                                                ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_36 (
                                                .CLKA(clka),      // Port A Clock
                                                .DOA(douta[36]),  // Port A 1-bit Data Output
                                                .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                .DIA(dina[36]),   // Port A 1-bit Data Input
                                                .ENA(ena[4]),    // Port A RAM Enable Input
                                                .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                .WEA(wea),         // Port A Write Enable Input
                                                .CLKB(clkb),      // Port B Clock
                                                .DOB(doutb[36]),  // Port B 1-bit Data Output
                                                .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                .DIB(dinb[36]),   // Port B 1-bit Data Input
                                                .ENB(enb[4]),    // Port B RAM Enable Input
                                                .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                .WEB(web)         // Port B Write Enable Input
                                                ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_37 (
                                                .CLKA(clka),      // Port A Clock
                                                .DOA(douta[37]),  // Port A 1-bit Data Output
                                                .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                .DIA(dina[37]),   // Port A 1-bit Data Input
                                                .ENA(ena[4]),    // Port A RAM Enable Input
                                                .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                .WEA(wea),         // Port A Write Enable Input
                                                .CLKB(clkb),      // Port B Clock
                                                .DOB(doutb[37]),  // Port B 1-bit Data Output
                                                .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                .DIB(dinb[37]),   // Port B 1-bit Data Input
                                                .ENB(enb[4]),    // Port B RAM Enable Input
                                                .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                .WEB(web)         // Port B Write Enable Input
                                                ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_38 (
                                                .CLKA(clka),      // Port A Clock
                                                .DOA(douta[38]),  // Port A 1-bit Data Output
                                                .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                .DIA(dina[38]),   // Port A 1-bit Data Input
                                                .ENA(ena[4]),    // Port A RAM Enable Input
                                                .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                .WEA(wea),         // Port A Write Enable Input
                                                .CLKB(clkb),      // Port B Clock
                                                .DOB(doutb[38]),  // Port B 1-bit Data Output
                                                .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                .DIB(dinb[38]),   // Port B 1-bit Data Input
                                                .ENB(enb[4]),    // Port B RAM Enable Input
                                                .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                .WEB(web)         // Port B Write Enable Input
                                                ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_39 (
                                                .CLKA(clka),      // Port A Clock
                                                .DOA(douta[39]),  // Port A 1-bit Data Output
                                                .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                .DIA(dina[39]),   // Port A 1-bit Data Input
                                                .ENA(ena[4]),    // Port A RAM Enable Input
                                                .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                .WEA(wea),         // Port A Write Enable Input
                                                .CLKB(clkb),      // Port B Clock
                                                .DOB(doutb[39]),  // Port B 1-bit Data Output
                                                .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                .DIB(dinb[39]),   // Port B 1-bit Data Input
                                                .ENB(enb[4]),    // Port B RAM Enable Input
                                                .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                .WEB(web)         // Port B Write Enable Input
                                                ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_40 (
                                                .CLKA(clka),      // Port A Clock
                                                .DOA(douta[40]),  // Port A 1-bit Data Output
                                                .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                .DIA(dina[40]),   // Port A 1-bit Data Input
                                                .ENA(ena[5]),    // Port A RAM Enable Input
                                                .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                .WEA(wea),         // Port A Write Enable Input
                                                .CLKB(clkb),      // Port B Clock
                                                .DOB(doutb[40]),  // Port B 1-bit Data Output
                                                .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                .DIB(dinb[40]),   // Port B 1-bit Data Input
                                                .ENB(enb[5]),    // Port B RAM Enable Input
                                                .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                .WEB(web)         // Port B Write Enable Input
                                                ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_41 (
                                                .CLKA(clka),      // Port A Clock
                                                .DOA(douta[41]),  // Port A 1-bit Data Output
                                                .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                .DIA(dina[41]),   // Port A 1-bit Data Input
                                                .ENA(ena[5]),    // Port A RAM Enable Input
                                                .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                .WEA(wea),         // Port A Write Enable Input
                                                .CLKB(clkb),      // Port B Clock
                                                .DOB(doutb[41]),  // Port B 1-bit Data Output
                                                .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                .DIB(dinb[41]),   // Port B 1-bit Data Input
                                                .ENB(enb[5]),    // Port B RAM Enable Input
                                                .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                .WEB(web)         // Port B Write Enable Input
                                                ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_42 (
                                                .CLKA(clka),      // Port A Clock
                                                .DOA(douta[42]),  // Port A 1-bit Data Output
                                                .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                .DIA(dina[42]),   // Port A 1-bit Data Input
                                                .ENA(ena[5]),    // Port A RAM Enable Input
                                                .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                .WEA(wea),         // Port A Write Enable Input
                                                .CLKB(clkb),      // Port B Clock
                                                .DOB(doutb[42]),  // Port B 1-bit Data Output
                                                .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                .DIB(dinb[42]),   // Port B 1-bit Data Input
                                                .ENB(enb[5]),    // Port B RAM Enable Input
                                                .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                .WEB(web)         // Port B Write Enable Input
                                                ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_43 (
                                                .CLKA(clka),      // Port A Clock
                                                .DOA(douta[43]),  // Port A 1-bit Data Output
                                                .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                .DIA(dina[43]),   // Port A 1-bit Data Input
                                                .ENA(ena[5]),    // Port A RAM Enable Input
                                                .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                .WEA(wea),         // Port A Write Enable Input
                                                .CLKB(clkb),      // Port B Clock
                                                .DOB(doutb[43]),  // Port B 1-bit Data Output
                                                .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                .DIB(dinb[43]),   // Port B 1-bit Data Input
                                                .ENB(enb[5]),    // Port B RAM Enable Input
                                                .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                .WEB(web)         // Port B Write Enable Input
                                                ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_44 (
                                                .CLKA(clka),      // Port A Clock
                                                .DOA(douta[44]),  // Port A 1-bit Data Output
                                                .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                .DIA(dina[44]),   // Port A 1-bit Data Input
                                                .ENA(ena[5]),    // Port A RAM Enable Input
                                                .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                .WEA(wea),         // Port A Write Enable Input
                                                .CLKB(clkb),      // Port B Clock
                                                .DOB(doutb[44]),  // Port B 1-bit Data Output
                                                .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                .DIB(dinb[44]),   // Port B 1-bit Data Input
                                                .ENB(enb[5]),    // Port B RAM Enable Input
                                                .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                .WEB(web)         // Port B Write Enable Input
                                                ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_45 (
                                                .CLKA(clka),      // Port A Clock
                                                .DOA(douta[45]),  // Port A 1-bit Data Output
                                                .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                .DIA(dina[45]),   // Port A 1-bit Data Input
                                                .ENA(ena[5]),    // Port A RAM Enable Input
                                                .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                .WEA(wea),         // Port A Write Enable Input
                                                .CLKB(clkb),      // Port B Clock
                                                .DOB(doutb[45]),  // Port B 1-bit Data Output
                                                .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                .DIB(dinb[45]),   // Port B 1-bit Data Input
                                                .ENB(enb[5]),    // Port B RAM Enable Input
                                                .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                .WEB(web)         // Port B Write Enable Input
                                                ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_46 (
                                                .CLKA(clka),      // Port A Clock
                                                .DOA(douta[46]),  // Port A 1-bit Data Output
                                                .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                .DIA(dina[46]),   // Port A 1-bit Data Input
                                                .ENA(ena[5]),    // Port A RAM Enable Input
                                                .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                .WEA(wea),         // Port A Write Enable Input
                                                .CLKB(clkb),      // Port B Clock
                                                .DOB(doutb[46]),  // Port B 1-bit Data Output
                                                .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                .DIB(dinb[46]),   // Port B 1-bit Data Input
                                                .ENB(enb[5]),    // Port B RAM Enable Input
                                                .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                .WEB(web)         // Port B Write Enable Input
                                                ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_47 (
                                                .CLKA(clka),      // Port A Clock
                                                .DOA(douta[47]),  // Port A 1-bit Data Output
                                                .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                .DIA(dina[47]),   // Port A 1-bit Data Input
                                                .ENA(ena[5]),    // Port A RAM Enable Input
                                                .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                .WEA(wea),         // Port A Write Enable Input
                                                .CLKB(clkb),      // Port B Clock
                                                .DOB(doutb[47]),  // Port B 1-bit Data Output
                                                .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                .DIB(dinb[47]),   // Port B 1-bit Data Input
                                                .ENB(enb[5]),    // Port B RAM Enable Input
                                                .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                .WEB(web)         // Port B Write Enable Input
                                                ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_48 (
                                                .CLKA(clka),      // Port A Clock
                                                .DOA(douta[48]),  // Port A 1-bit Data Output
                                                .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                .DIA(dina[48]),   // Port A 1-bit Data Input
                                                .ENA(ena[6]),    // Port A RAM Enable Input
                                                .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                .WEA(wea),         // Port A Write Enable Input
                                                .CLKB(clkb),      // Port B Clock
                                                .DOB(doutb[48]),  // Port B 1-bit Data Output
                                                .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                .DIB(dinb[48]),   // Port B 1-bit Data Input
                                                .ENB(enb[6]),    // Port B RAM Enable Input
                                                .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                .WEB(web)         // Port B Write Enable Input
                                                ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_49 (
                                                .CLKA(clka),      // Port A Clock
                                                .DOA(douta[49]),  // Port A 1-bit Data Output
                                                .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                .DIA(dina[49]),   // Port A 1-bit Data Input
                                                .ENA(ena[6]),    // Port A RAM Enable Input
                                                .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                .WEA(wea),         // Port A Write Enable Input
                                                .CLKB(clkb),      // Port B Clock
                                                .DOB(doutb[49]),  // Port B 1-bit Data Output
                                                .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                .DIB(dinb[49]),   // Port B 1-bit Data Input
                                                .ENB(enb[6]),    // Port B RAM Enable Input
                                                .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                .WEB(web)         // Port B Write Enable Input
                                                ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_50 (
                                                .CLKA(clka),      // Port A Clock
                                                .DOA(douta[50]),  // Port A 1-bit Data Output
                                                .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                .DIA(dina[50]),   // Port A 1-bit Data Input
                                                .ENA(ena[6]),    // Port A RAM Enable Input
                                                .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                .WEA(wea),         // Port A Write Enable Input
                                                .CLKB(clkb),      // Port B Clock
                                                .DOB(doutb[50]),  // Port B 1-bit Data Output
                                                .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                .DIB(dinb[50]),   // Port B 1-bit Data Input
                                                .ENB(enb[6]),    // Port B RAM Enable Input
                                                .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                .WEB(web)         // Port B Write Enable Input
                                                ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_51 (
                                                .CLKA(clka),      // Port A Clock
                                                .DOA(douta[51]),  // Port A 1-bit Data Output
                                                .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                .DIA(dina[51]),   // Port A 1-bit Data Input
                                                .ENA(ena[6]),    // Port A RAM Enable Input
                                                .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                .WEA(wea),         // Port A Write Enable Input
                                                .CLKB(clkb),      // Port B Clock
                                                .DOB(doutb[51]),  // Port B 1-bit Data Output
                                                .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                .DIB(dinb[51]),   // Port B 1-bit Data Input
                                                .ENB(enb[6]),    // Port B RAM Enable Input
                                                .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                .WEB(web)         // Port B Write Enable Input
                                                ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_52 (
                                                .CLKA(clka),      // Port A Clock
                                                .DOA(douta[52]),  // Port A 1-bit Data Output
                                                .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                .DIA(dina[52]),   // Port A 1-bit Data Input
                                                .ENA(ena[6]),    // Port A RAM Enable Input
                                                .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                .WEA(wea),         // Port A Write Enable Input
                                                .CLKB(clkb),      // Port B Clock
                                                .DOB(doutb[52]),  // Port B 1-bit Data Output
                                                .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                .DIB(dinb[52]),   // Port B 1-bit Data Input
                                                .ENB(enb[6]),    // Port B RAM Enable Input
                                                .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                .WEB(web)         // Port B Write Enable Input
                                                ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_53 (
                                                .CLKA(clka),      // Port A Clock
                                                .DOA(douta[53]),  // Port A 1-bit Data Output
                                                .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                .DIA(dina[53]),   // Port A 1-bit Data Input
                                                .ENA(ena[6]),    // Port A RAM Enable Input
                                                .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                .WEA(wea),         // Port A Write Enable Input
                                                .CLKB(clkb),      // Port B Clock
                                                .DOB(doutb[53]),  // Port B 1-bit Data Output
                                                .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                .DIB(dinb[53]),   // Port B 1-bit Data Input
                                                .ENB(enb[6]),    // Port B RAM Enable Input
                                                .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                .WEB(web)         // Port B Write Enable Input
                                                ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_54 (
                                                .CLKA(clka),      // Port A Clock
                                                .DOA(douta[54]),  // Port A 1-bit Data Output
                                                .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                .DIA(dina[54]),   // Port A 1-bit Data Input
                                                .ENA(ena[6]),    // Port A RAM Enable Input
                                                .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                .WEA(wea),         // Port A Write Enable Input
                                                .CLKB(clkb),      // Port B Clock
                                                .DOB(doutb[54]),  // Port B 1-bit Data Output
                                                .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                .DIB(dinb[54]),   // Port B 1-bit Data Input
                                                .ENB(enb[6]),    // Port B RAM Enable Input
                                                .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                .WEB(web)         // Port B Write Enable Input
                                                ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_55 (
                                                .CLKA(clka),      // Port A Clock
                                                .DOA(douta[55]),  // Port A 1-bit Data Output
                                                .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                .DIA(dina[55]),   // Port A 1-bit Data Input
                                                .ENA(ena[6]),    // Port A RAM Enable Input
                                                .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                .WEA(wea),         // Port A Write Enable Input
                                                .CLKB(clkb),      // Port B Clock
                                                .DOB(doutb[55]),  // Port B 1-bit Data Output
                                                .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                .DIB(dinb[55]),   // Port B 1-bit Data Input
                                                .ENB(enb[6]),    // Port B RAM Enable Input
                                                .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                .WEB(web)         // Port B Write Enable Input
                                                ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_56 (
                                                .CLKA(clka),      // Port A Clock
                                                .DOA(douta[56]),  // Port A 1-bit Data Output
                                                .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                .DIA(dina[56]),   // Port A 1-bit Data Input
                                                .ENA(ena[7]),    // Port A RAM Enable Input
                                                .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                .WEA(wea),         // Port A Write Enable Input
                                                .CLKB(clkb),      // Port B Clock
                                                .DOB(doutb[56]),  // Port B 1-bit Data Output
                                                .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                .DIB(dinb[56]),   // Port B 1-bit Data Input
                                                .ENB(enb[7]),    // Port B RAM Enable Input
                                                .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                .WEB(web)         // Port B Write Enable Input
                                                ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_57 (
                                                .CLKA(clka),      // Port A Clock
                                                .DOA(douta[57]),  // Port A 1-bit Data Output
                                                .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                .DIA(dina[57]),   // Port A 1-bit Data Input
                                                .ENA(ena[7]),    // Port A RAM Enable Input
                                                .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                .WEA(wea),         // Port A Write Enable Input
                                                .CLKB(clkb),      // Port B Clock
                                                .DOB(doutb[57]),  // Port B 1-bit Data Output
                                                .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                .DIB(dinb[57]),   // Port B 1-bit Data Input
                                                .ENB(enb[7]),    // Port B RAM Enable Input
                                                .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                .WEB(web)         // Port B Write Enable Input
                                                ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_58 (
                                                .CLKA(clka),      // Port A Clock
                                                .DOA(douta[58]),  // Port A 1-bit Data Output
                                                .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                .DIA(dina[58]),   // Port A 1-bit Data Input
                                                .ENA(ena[7]),    // Port A RAM Enable Input
                                                .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                .WEA(wea),         // Port A Write Enable Input
                                                .CLKB(clkb),      // Port B Clock
                                                .DOB(doutb[58]),  // Port B 1-bit Data Output
                                                .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                .DIB(dinb[58]),   // Port B 1-bit Data Input
                                                .ENB(enb[7]),    // Port B RAM Enable Input
                                                .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                .WEB(web)         // Port B Write Enable Input
                                                ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_59 (
                                                .CLKA(clka),      // Port A Clock
                                                .DOA(douta[59]),  // Port A 1-bit Data Output
                                                .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                .DIA(dina[59]),   // Port A 1-bit Data Input
                                                .ENA(ena[7]),    // Port A RAM Enable Input
                                                .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                .WEA(wea),         // Port A Write Enable Input
                                                .CLKB(clkb),      // Port B Clock
                                                .DOB(doutb[59]),  // Port B 1-bit Data Output
                                                .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                .DIB(dinb[59]),   // Port B 1-bit Data Input
                                                .ENB(enb[7]),    // Port B RAM Enable Input
                                                .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                .WEB(web)         // Port B Write Enable Input
                                                ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_60 (
                                                .CLKA(clka),      // Port A Clock
                                                .DOA(douta[60]),  // Port A 1-bit Data Output
                                                .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                .DIA(dina[60]),   // Port A 1-bit Data Input
                                                .ENA(ena[7]),    // Port A RAM Enable Input
                                                .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                .WEA(wea),         // Port A Write Enable Input
                                                .CLKB(clkb),      // Port B Clock
                                                .DOB(doutb[60]),  // Port B 1-bit Data Output
                                                .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                .DIB(dinb[60]),   // Port B 1-bit Data Input
                                                .ENB(enb[7]),    // Port B RAM Enable Input
                                                .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                .WEB(web)         // Port B Write Enable Input
                                                ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_61 (
                                                .CLKA(clka),      // Port A Clock
                                                .DOA(douta[61]),  // Port A 1-bit Data Output
                                                .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                .DIA(dina[61]),   // Port A 1-bit Data Input
                                                .ENA(ena[7]),    // Port A RAM Enable Input
                                                .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                .WEA(wea),         // Port A Write Enable Input
                                                .CLKB(clkb),      // Port B Clock
                                                .DOB(doutb[61]),  // Port B 1-bit Data Output
                                                .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                .DIB(dinb[61]),   // Port B 1-bit Data Input
                                                .ENB(enb[7]),    // Port B RAM Enable Input
                                                .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                .WEB(web)         // Port B Write Enable Input
                                                ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_62 (
                                                .CLKA(clka),      // Port A Clock
                                                .DOA(douta[62]),  // Port A 1-bit Data Output
                                                .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                .DIA(dina[62]),   // Port A 1-bit Data Input
                                                .ENA(ena[7]),    // Port A RAM Enable Input
                                                .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                .WEA(wea),         // Port A Write Enable Input
                                                .CLKB(clkb),      // Port B Clock
                                                .DOB(doutb[62]),  // Port B 1-bit Data Output
                                                .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                .DIB(dinb[62]),   // Port B 1-bit Data Input
                                                .ENB(enb[7]),    // Port B RAM Enable Input
                                                .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                .WEB(web)         // Port B Write Enable Input
                                                ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_63 (
                                                .CLKA(clka),      // Port A Clock
                                                .DOA(douta[63]),  // Port A 1-bit Data Output
                                                .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                .DIA(dina[63]),   // Port A 1-bit Data Input
                                                .ENA(ena[7]),    // Port A RAM Enable Input
                                                .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                .WEA(wea),         // Port A Write Enable Input
                                                .CLKB(clkb),      // Port B Clock
                                                .DOB(doutb[63]),  // Port B 1-bit Data Output
                                                .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                .DIB(dinb[63]),   // Port B 1-bit Data Input
                                                .ENB(enb[7]),    // Port B RAM Enable Input
                                                .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                .WEB(web)         // Port B Write Enable Input
                                                ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_64 (
                                                .CLKA(clka),      // Port A Clock
                                                .DOA(douta[64]),  // Port A 1-bit Data Output
                                                .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                .DIA(dina[64]),   // Port A 1-bit Data Input
                                                .ENA(ena[8]),    // Port A RAM Enable Input
                                                .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                .WEA(wea),         // Port A Write Enable Input
                                                .CLKB(clkb),      // Port B Clock
                                                .DOB(doutb[64]),  // Port B 1-bit Data Output
                                                .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                .DIB(dinb[64]),   // Port B 1-bit Data Input
                                                .ENB(enb[8]),    // Port B RAM Enable Input
                                                .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                .WEB(web)         // Port B Write Enable Input
                                                ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_65 (
                                                .CLKA(clka),      // Port A Clock
                                                .DOA(douta[65]),  // Port A 1-bit Data Output
                                                .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                .DIA(dina[65]),   // Port A 1-bit Data Input
                                                .ENA(ena[8]),    // Port A RAM Enable Input
                                                .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                .WEA(wea),         // Port A Write Enable Input
                                                .CLKB(clkb),      // Port B Clock
                                                .DOB(doutb[65]),  // Port B 1-bit Data Output
                                                .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                .DIB(dinb[65]),   // Port B 1-bit Data Input
                                                .ENB(enb[8]),    // Port B RAM Enable Input
                                                .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                .WEB(web)         // Port B Write Enable Input
                                                ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_66 (
                                                .CLKA(clka),      // Port A Clock
                                                .DOA(douta[66]),  // Port A 1-bit Data Output
                                                .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                .DIA(dina[66]),   // Port A 1-bit Data Input
                                                .ENA(ena[8]),    // Port A RAM Enable Input
                                                .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                .WEA(wea),         // Port A Write Enable Input
                                                .CLKB(clkb),      // Port B Clock
                                                .DOB(doutb[66]),  // Port B 1-bit Data Output
                                                .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                .DIB(dinb[66]),   // Port B 1-bit Data Input
                                                .ENB(enb[8]),    // Port B RAM Enable Input
                                                .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                .WEB(web)         // Port B Write Enable Input
                                                ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_67 (
                                                .CLKA(clka),      // Port A Clock
                                                .DOA(douta[67]),  // Port A 1-bit Data Output
                                                .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                .DIA(dina[67]),   // Port A 1-bit Data Input
                                                .ENA(ena[8]),    // Port A RAM Enable Input
                                                .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                .WEA(wea),         // Port A Write Enable Input
                                                .CLKB(clkb),      // Port B Clock
                                                .DOB(doutb[67]),  // Port B 1-bit Data Output
                                                .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                .DIB(dinb[67]),   // Port B 1-bit Data Input
                                                .ENB(enb[8]),    // Port B RAM Enable Input
                                                .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                .WEB(web)         // Port B Write Enable Input
                                                ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_68 (
                                                .CLKA(clka),      // Port A Clock
                                                .DOA(douta[68]),  // Port A 1-bit Data Output
                                                .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                .DIA(dina[68]),   // Port A 1-bit Data Input
                                                .ENA(ena[8]),    // Port A RAM Enable Input
                                                .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                .WEA(wea),         // Port A Write Enable Input
                                                .CLKB(clkb),      // Port B Clock
                                                .DOB(doutb[68]),  // Port B 1-bit Data Output
                                                .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                .DIB(dinb[68]),   // Port B 1-bit Data Input
                                                .ENB(enb[8]),    // Port B RAM Enable Input
                                                .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                .WEB(web)         // Port B Write Enable Input
                                                ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_69 (
                                                .CLKA(clka),      // Port A Clock
                                                .DOA(douta[69]),  // Port A 1-bit Data Output
                                                .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                .DIA(dina[69]),   // Port A 1-bit Data Input
                                                .ENA(ena[8]),    // Port A RAM Enable Input
                                                .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                .WEA(wea),         // Port A Write Enable Input
                                                .CLKB(clkb),      // Port B Clock
                                                .DOB(doutb[69]),  // Port B 1-bit Data Output
                                                .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                .DIB(dinb[69]),   // Port B 1-bit Data Input
                                                .ENB(enb[8]),    // Port B RAM Enable Input
                                                .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                .WEB(web)         // Port B Write Enable Input
                                                ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_70 (
                                                .CLKA(clka),      // Port A Clock
                                                .DOA(douta[70]),  // Port A 1-bit Data Output
                                                .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                .DIA(dina[70]),   // Port A 1-bit Data Input
                                                .ENA(ena[8]),    // Port A RAM Enable Input
                                                .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                .WEA(wea),         // Port A Write Enable Input
                                                .CLKB(clkb),      // Port B Clock
                                                .DOB(doutb[70]),  // Port B 1-bit Data Output
                                                .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                .DIB(dinb[70]),   // Port B 1-bit Data Input
                                                .ENB(enb[8]),    // Port B RAM Enable Input
                                                .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                .WEB(web)         // Port B Write Enable Input
                                                ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_71 (
                                                .CLKA(clka),      // Port A Clock
                                                .DOA(douta[71]),  // Port A 1-bit Data Output
                                                .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                .DIA(dina[71]),   // Port A 1-bit Data Input
                                                .ENA(ena[8]),    // Port A RAM Enable Input
                                                .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                .WEA(wea),         // Port A Write Enable Input
                                                .CLKB(clkb),      // Port B Clock
                                                .DOB(doutb[71]),  // Port B 1-bit Data Output
                                                .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                .DIB(dinb[71]),   // Port B 1-bit Data Input
                                                .ENB(enb[8]),    // Port B RAM Enable Input
                                                .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                .WEB(web)         // Port B Write Enable Input
                                                ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_72 (
                                                .CLKA(clka),      // Port A Clock
                                                .DOA(douta[72]),  // Port A 1-bit Data Output
                                                .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                .DIA(dina[72]),   // Port A 1-bit Data Input
                                                .ENA(ena[9]),    // Port A RAM Enable Input
                                                .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                .WEA(wea),         // Port A Write Enable Input
                                                .CLKB(clkb),      // Port B Clock
                                                .DOB(doutb[72]),  // Port B 1-bit Data Output
                                                .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                .DIB(dinb[72]),   // Port B 1-bit Data Input
                                                .ENB(enb[9]),    // Port B RAM Enable Input
                                                .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                .WEB(web)         // Port B Write Enable Input
                                                ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_73 (
                                                .CLKA(clka),      // Port A Clock
                                                .DOA(douta[73]),  // Port A 1-bit Data Output
                                                .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                .DIA(dina[73]),   // Port A 1-bit Data Input
                                                .ENA(ena[9]),    // Port A RAM Enable Input
                                                .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                .WEA(wea),         // Port A Write Enable Input
                                                .CLKB(clkb),      // Port B Clock
                                                .DOB(doutb[73]),  // Port B 1-bit Data Output
                                                .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                .DIB(dinb[73]),   // Port B 1-bit Data Input
                                                .ENB(enb[9]),    // Port B RAM Enable Input
                                                .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                .WEB(web)         // Port B Write Enable Input
                                                ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_74 (
                                                .CLKA(clka),      // Port A Clock
                                                .DOA(douta[74]),  // Port A 1-bit Data Output
                                                .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                .DIA(dina[74]),   // Port A 1-bit Data Input
                                                .ENA(ena[9]),    // Port A RAM Enable Input
                                                .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                .WEA(wea),         // Port A Write Enable Input
                                                .CLKB(clkb),      // Port B Clock
                                                .DOB(doutb[74]),  // Port B 1-bit Data Output
                                                .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                .DIB(dinb[74]),   // Port B 1-bit Data Input
                                                .ENB(enb[9]),    // Port B RAM Enable Input
                                                .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                .WEB(web)         // Port B Write Enable Input
                                                ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_75 (
                                                .CLKA(clka),      // Port A Clock
                                                .DOA(douta[75]),  // Port A 1-bit Data Output
                                                .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                .DIA(dina[75]),   // Port A 1-bit Data Input
                                                .ENA(ena[9]),    // Port A RAM Enable Input
                                                .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                .WEA(wea),         // Port A Write Enable Input
                                                .CLKB(clkb),      // Port B Clock
                                                .DOB(doutb[75]),  // Port B 1-bit Data Output
                                                .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                .DIB(dinb[75]),   // Port B 1-bit Data Input
                                                .ENB(enb[9]),    // Port B RAM Enable Input
                                                .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                .WEB(web)         // Port B Write Enable Input
                                                ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_76 (
                                                .CLKA(clka),      // Port A Clock
                                                .DOA(douta[76]),  // Port A 1-bit Data Output
                                                .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                .DIA(dina[76]),   // Port A 1-bit Data Input
                                                .ENA(ena[9]),    // Port A RAM Enable Input
                                                .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                .WEA(wea),         // Port A Write Enable Input
                                                .CLKB(clkb),      // Port B Clock
                                                .DOB(doutb[76]),  // Port B 1-bit Data Output
                                                .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                .DIB(dinb[76]),   // Port B 1-bit Data Input
                                                .ENB(enb[9]),    // Port B RAM Enable Input
                                                .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                .WEB(web)         // Port B Write Enable Input
                                                ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_77 (
                                                .CLKA(clka),      // Port A Clock
                                                .DOA(douta[77]),  // Port A 1-bit Data Output
                                                .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                .DIA(dina[77]),   // Port A 1-bit Data Input
                                                .ENA(ena[9]),    // Port A RAM Enable Input
                                                .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                .WEA(wea),         // Port A Write Enable Input
                                                .CLKB(clkb),      // Port B Clock
                                                .DOB(doutb[77]),  // Port B 1-bit Data Output
                                                .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                .DIB(dinb[77]),   // Port B 1-bit Data Input
                                                .ENB(enb[9]),    // Port B RAM Enable Input
                                                .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                .WEB(web)         // Port B Write Enable Input
                                                ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_78 (
                                                .CLKA(clka),      // Port A Clock
                                                .DOA(douta[78]),  // Port A 1-bit Data Output
                                                .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                .DIA(dina[78]),   // Port A 1-bit Data Input
                                                .ENA(ena[9]),    // Port A RAM Enable Input
                                                .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                .WEA(wea),         // Port A Write Enable Input
                                                .CLKB(clkb),      // Port B Clock
                                                .DOB(doutb[78]),  // Port B 1-bit Data Output
                                                .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                .DIB(dinb[78]),   // Port B 1-bit Data Input
                                                .ENB(enb[9]),    // Port B RAM Enable Input
                                                .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                .WEB(web)         // Port B Write Enable Input
                                                ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_79 (
                                                .CLKA(clka),      // Port A Clock
                                                .DOA(douta[79]),  // Port A 1-bit Data Output
                                                .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                .DIA(dina[79]),   // Port A 1-bit Data Input
                                                .ENA(ena[9]),    // Port A RAM Enable Input
                                                .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                .WEA(wea),         // Port A Write Enable Input
                                                .CLKB(clkb),      // Port B Clock
                                                .DOB(doutb[79]),  // Port B 1-bit Data Output
                                                .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                .DIB(dinb[79]),   // Port B 1-bit Data Input
                                                .ENB(enb[9]),    // Port B RAM Enable Input
                                                .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                .WEB(web)         // Port B Write Enable Input
                                                ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_80 (
                                                .CLKA(clka),      // Port A Clock
                                                .DOA(douta[80]),  // Port A 1-bit Data Output
                                                .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                .DIA(dina[80]),   // Port A 1-bit Data Input
                                                .ENA(ena[10]),    // Port A RAM Enable Input
                                                .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                .WEA(wea),         // Port A Write Enable Input
                                                .CLKB(clkb),      // Port B Clock
                                                .DOB(doutb[80]),  // Port B 1-bit Data Output
                                                .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                .DIB(dinb[80]),   // Port B 1-bit Data Input
                                                .ENB(enb[10]),    // Port B RAM Enable Input
                                                .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                .WEB(web)         // Port B Write Enable Input
                                                ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_81 (
                                                .CLKA(clka),      // Port A Clock
                                                .DOA(douta[81]),  // Port A 1-bit Data Output
                                                .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                .DIA(dina[81]),   // Port A 1-bit Data Input
                                                .ENA(ena[10]),    // Port A RAM Enable Input
                                                .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                .WEA(wea),         // Port A Write Enable Input
                                                .CLKB(clkb),      // Port B Clock
                                                .DOB(doutb[81]),  // Port B 1-bit Data Output
                                                .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                .DIB(dinb[81]),   // Port B 1-bit Data Input
                                                .ENB(enb[10]),    // Port B RAM Enable Input
                                                .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                .WEB(web)         // Port B Write Enable Input
                                                ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_82 (
                                                .CLKA(clka),      // Port A Clock
                                                .DOA(douta[82]),  // Port A 1-bit Data Output
                                                .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                .DIA(dina[82]),   // Port A 1-bit Data Input
                                                .ENA(ena[10]),    // Port A RAM Enable Input
                                                .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                .WEA(wea),         // Port A Write Enable Input
                                                .CLKB(clkb),      // Port B Clock
                                                .DOB(doutb[82]),  // Port B 1-bit Data Output
                                                .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                .DIB(dinb[82]),   // Port B 1-bit Data Input
                                                .ENB(enb[10]),    // Port B RAM Enable Input
                                                .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                .WEB(web)         // Port B Write Enable Input
                                                ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_83 (
                                                .CLKA(clka),      // Port A Clock
                                                .DOA(douta[83]),  // Port A 1-bit Data Output
                                                .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                .DIA(dina[83]),   // Port A 1-bit Data Input
                                                .ENA(ena[10]),    // Port A RAM Enable Input
                                                .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                .WEA(wea),         // Port A Write Enable Input
                                                .CLKB(clkb),      // Port B Clock
                                                .DOB(doutb[83]),  // Port B 1-bit Data Output
                                                .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                .DIB(dinb[83]),   // Port B 1-bit Data Input
                                                .ENB(enb[10]),    // Port B RAM Enable Input
                                                .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                .WEB(web)         // Port B Write Enable Input
                                                ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_84 (
                                                .CLKA(clka),      // Port A Clock
                                                .DOA(douta[84]),  // Port A 1-bit Data Output
                                                .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                .DIA(dina[84]),   // Port A 1-bit Data Input
                                                .ENA(ena[10]),    // Port A RAM Enable Input
                                                .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                .WEA(wea),         // Port A Write Enable Input
                                                .CLKB(clkb),      // Port B Clock
                                                .DOB(doutb[84]),  // Port B 1-bit Data Output
                                                .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                .DIB(dinb[84]),   // Port B 1-bit Data Input
                                                .ENB(enb[10]),    // Port B RAM Enable Input
                                                .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                .WEB(web)         // Port B Write Enable Input
                                                ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_85 (
                                                .CLKA(clka),      // Port A Clock
                                                .DOA(douta[85]),  // Port A 1-bit Data Output
                                                .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                .DIA(dina[85]),   // Port A 1-bit Data Input
                                                .ENA(ena[10]),    // Port A RAM Enable Input
                                                .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                .WEA(wea),         // Port A Write Enable Input
                                                .CLKB(clkb),      // Port B Clock
                                                .DOB(doutb[85]),  // Port B 1-bit Data Output
                                                .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                .DIB(dinb[85]),   // Port B 1-bit Data Input
                                                .ENB(enb[10]),    // Port B RAM Enable Input
                                                .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                .WEB(web)         // Port B Write Enable Input
                                                ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_86 (
                                                .CLKA(clka),      // Port A Clock
                                                .DOA(douta[86]),  // Port A 1-bit Data Output
                                                .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                .DIA(dina[86]),   // Port A 1-bit Data Input
                                                .ENA(ena[10]),    // Port A RAM Enable Input
                                                .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                .WEA(wea),         // Port A Write Enable Input
                                                .CLKB(clkb),      // Port B Clock
                                                .DOB(doutb[86]),  // Port B 1-bit Data Output
                                                .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                .DIB(dinb[86]),   // Port B 1-bit Data Input
                                                .ENB(enb[10]),    // Port B RAM Enable Input
                                                .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                .WEB(web)         // Port B Write Enable Input
                                                ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_87 (
                                                .CLKA(clka),      // Port A Clock
                                                .DOA(douta[87]),  // Port A 1-bit Data Output
                                                .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                .DIA(dina[87]),   // Port A 1-bit Data Input
                                                .ENA(ena[10]),    // Port A RAM Enable Input
                                                .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                .WEA(wea),         // Port A Write Enable Input
                                                .CLKB(clkb),      // Port B Clock
                                                .DOB(doutb[87]),  // Port B 1-bit Data Output
                                                .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                .DIB(dinb[87]),   // Port B 1-bit Data Input
                                                .ENB(enb[10]),    // Port B RAM Enable Input
                                                .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                .WEB(web)         // Port B Write Enable Input
                                                ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_88 (
                                                .CLKA(clka),      // Port A Clock
                                                .DOA(douta[88]),  // Port A 1-bit Data Output
                                                .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                .DIA(dina[88]),   // Port A 1-bit Data Input
                                                .ENA(ena[11]),    // Port A RAM Enable Input
                                                .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                .WEA(wea),         // Port A Write Enable Input
                                                .CLKB(clkb),      // Port B Clock
                                                .DOB(doutb[88]),  // Port B 1-bit Data Output
                                                .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                .DIB(dinb[88]),   // Port B 1-bit Data Input
                                                .ENB(enb[11]),    // Port B RAM Enable Input
                                                .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                .WEB(web)         // Port B Write Enable Input
                                                ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_89 (
                                                .CLKA(clka),      // Port A Clock
                                                .DOA(douta[89]),  // Port A 1-bit Data Output
                                                .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                .DIA(dina[89]),   // Port A 1-bit Data Input
                                                .ENA(ena[11]),    // Port A RAM Enable Input
                                                .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                .WEA(wea),         // Port A Write Enable Input
                                                .CLKB(clkb),      // Port B Clock
                                                .DOB(doutb[89]),  // Port B 1-bit Data Output
                                                .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                .DIB(dinb[89]),   // Port B 1-bit Data Input
                                                .ENB(enb[11]),    // Port B RAM Enable Input
                                                .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                .WEB(web)         // Port B Write Enable Input
                                                ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_90 (
                                                .CLKA(clka),      // Port A Clock
                                                .DOA(douta[90]),  // Port A 1-bit Data Output
                                                .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                .DIA(dina[90]),   // Port A 1-bit Data Input
                                                .ENA(ena[11]),    // Port A RAM Enable Input
                                                .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                .WEA(wea),         // Port A Write Enable Input
                                                .CLKB(clkb),      // Port B Clock
                                                .DOB(doutb[90]),  // Port B 1-bit Data Output
                                                .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                .DIB(dinb[90]),   // Port B 1-bit Data Input
                                                .ENB(enb[11]),    // Port B RAM Enable Input
                                                .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                .WEB(web)         // Port B Write Enable Input
                                                ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_91 (
                                                .CLKA(clka),      // Port A Clock
                                                .DOA(douta[91]),  // Port A 1-bit Data Output
                                                .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                .DIA(dina[91]),   // Port A 1-bit Data Input
                                                .ENA(ena[11]),    // Port A RAM Enable Input
                                                .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                .WEA(wea),         // Port A Write Enable Input
                                                .CLKB(clkb),      // Port B Clock
                                                .DOB(doutb[91]),  // Port B 1-bit Data Output
                                                .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                .DIB(dinb[91]),   // Port B 1-bit Data Input
                                                .ENB(enb[11]),    // Port B RAM Enable Input
                                                .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                .WEB(web)         // Port B Write Enable Input
                                                ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_92 (
                                                .CLKA(clka),      // Port A Clock
                                                .DOA(douta[92]),  // Port A 1-bit Data Output
                                                .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                .DIA(dina[92]),   // Port A 1-bit Data Input
                                                .ENA(ena[11]),    // Port A RAM Enable Input
                                                .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                .WEA(wea),         // Port A Write Enable Input
                                                .CLKB(clkb),      // Port B Clock
                                                .DOB(doutb[92]),  // Port B 1-bit Data Output
                                                .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                .DIB(dinb[92]),   // Port B 1-bit Data Input
                                                .ENB(enb[11]),    // Port B RAM Enable Input
                                                .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                .WEB(web)         // Port B Write Enable Input
                                                ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_93 (
                                                .CLKA(clka),      // Port A Clock
                                                .DOA(douta[93]),  // Port A 1-bit Data Output
                                                .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                .DIA(dina[93]),   // Port A 1-bit Data Input
                                                .ENA(ena[11]),    // Port A RAM Enable Input
                                                .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                .WEA(wea),         // Port A Write Enable Input
                                                .CLKB(clkb),      // Port B Clock
                                                .DOB(doutb[93]),  // Port B 1-bit Data Output
                                                .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                .DIB(dinb[93]),   // Port B 1-bit Data Input
                                                .ENB(enb[11]),    // Port B RAM Enable Input
                                                .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                .WEB(web)         // Port B Write Enable Input
                                                ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_94 (
                                                .CLKA(clka),      // Port A Clock
                                                .DOA(douta[94]),  // Port A 1-bit Data Output
                                                .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                .DIA(dina[94]),   // Port A 1-bit Data Input
                                                .ENA(ena[11]),    // Port A RAM Enable Input
                                                .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                .WEA(wea),         // Port A Write Enable Input
                                                .CLKB(clkb),      // Port B Clock
                                                .DOB(doutb[94]),  // Port B 1-bit Data Output
                                                .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                .DIB(dinb[94]),   // Port B 1-bit Data Input
                                                .ENB(enb[11]),    // Port B RAM Enable Input
                                                .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                .WEB(web)         // Port B Write Enable Input
                                                ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_95 (
                                                .CLKA(clka),      // Port A Clock
                                                .DOA(douta[95]),  // Port A 1-bit Data Output
                                                .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                .DIA(dina[95]),   // Port A 1-bit Data Input
                                                .ENA(ena[11]),    // Port A RAM Enable Input
                                                .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                .WEA(wea),         // Port A Write Enable Input
                                                .CLKB(clkb),      // Port B Clock
                                                .DOB(doutb[95]),  // Port B 1-bit Data Output
                                                .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                .DIB(dinb[95]),   // Port B 1-bit Data Input
                                                .ENB(enb[11]),    // Port B RAM Enable Input
                                                .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                .WEB(web)         // Port B Write Enable Input
                                                ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_96 (
                                                .CLKA(clka),      // Port A Clock
                                                .DOA(douta[96]),  // Port A 1-bit Data Output
                                                .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                .DIA(dina[96]),   // Port A 1-bit Data Input
                                                .ENA(ena[12]),    // Port A RAM Enable Input
                                                .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                .WEA(wea),         // Port A Write Enable Input
                                                .CLKB(clkb),      // Port B Clock
                                                .DOB(doutb[96]),  // Port B 1-bit Data Output
                                                .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                .DIB(dinb[96]),   // Port B 1-bit Data Input
                                                .ENB(enb[12]),    // Port B RAM Enable Input
                                                .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                .WEB(web)         // Port B Write Enable Input
                                                ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_97 (
                                                .CLKA(clka),      // Port A Clock
                                                .DOA(douta[97]),  // Port A 1-bit Data Output
                                                .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                .DIA(dina[97]),   // Port A 1-bit Data Input
                                                .ENA(ena[12]),    // Port A RAM Enable Input
                                                .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                .WEA(wea),         // Port A Write Enable Input
                                                .CLKB(clkb),      // Port B Clock
                                                .DOB(doutb[97]),  // Port B 1-bit Data Output
                                                .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                .DIB(dinb[97]),   // Port B 1-bit Data Input
                                                .ENB(enb[12]),    // Port B RAM Enable Input
                                                .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                .WEB(web)         // Port B Write Enable Input
                                                ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_98 (
                                                .CLKA(clka),      // Port A Clock
                                                .DOA(douta[98]),  // Port A 1-bit Data Output
                                                .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                .DIA(dina[98]),   // Port A 1-bit Data Input
                                                .ENA(ena[12]),    // Port A RAM Enable Input
                                                .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                .WEA(wea),         // Port A Write Enable Input
                                                .CLKB(clkb),      // Port B Clock
                                                .DOB(doutb[98]),  // Port B 1-bit Data Output
                                                .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                .DIB(dinb[98]),   // Port B 1-bit Data Input
                                                .ENB(enb[12]),    // Port B RAM Enable Input
                                                .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                .WEB(web)         // Port B Write Enable Input
                                                ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_99 (
                                                .CLKA(clka),      // Port A Clock
                                                .DOA(douta[99]),  // Port A 1-bit Data Output
                                                .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                .DIA(dina[99]),   // Port A 1-bit Data Input
                                                .ENA(ena[12]),    // Port A RAM Enable Input
                                                .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                .WEA(wea),         // Port A Write Enable Input
                                                .CLKB(clkb),      // Port B Clock
                                                .DOB(doutb[99]),  // Port B 1-bit Data Output
                                                .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                .DIB(dinb[99]),   // Port B 1-bit Data Input
                                                .ENB(enb[12]),    // Port B RAM Enable Input
                                                .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                .WEB(web)         // Port B Write Enable Input
                                                ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_100 (
                                                 .CLKA(clka),      // Port A Clock
                                                 .DOA(douta[100]),  // Port A 1-bit Data Output
                                                 .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                 .DIA(dina[100]),   // Port A 1-bit Data Input
                                                 .ENA(ena[12]),    // Port A RAM Enable Input
                                                 .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                 .WEA(wea),         // Port A Write Enable Input
                                                 .CLKB(clkb),      // Port B Clock
                                                 .DOB(doutb[100]),  // Port B 1-bit Data Output
                                                 .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                 .DIB(dinb[100]),   // Port B 1-bit Data Input
                                                 .ENB(enb[12]),    // Port B RAM Enable Input
                                                 .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                 .WEB(web)         // Port B Write Enable Input
                                                 ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_101 (
                                                 .CLKA(clka),      // Port A Clock
                                                 .DOA(douta[101]),  // Port A 1-bit Data Output
                                                 .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                 .DIA(dina[101]),   // Port A 1-bit Data Input
                                                 .ENA(ena[12]),    // Port A RAM Enable Input
                                                 .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                 .WEA(wea),         // Port A Write Enable Input
                                                 .CLKB(clkb),      // Port B Clock
                                                 .DOB(doutb[101]),  // Port B 1-bit Data Output
                                                 .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                 .DIB(dinb[101]),   // Port B 1-bit Data Input
                                                 .ENB(enb[12]),    // Port B RAM Enable Input
                                                 .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                 .WEB(web)         // Port B Write Enable Input
                                                 ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_102 (
                                                 .CLKA(clka),      // Port A Clock
                                                 .DOA(douta[102]),  // Port A 1-bit Data Output
                                                 .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                 .DIA(dina[102]),   // Port A 1-bit Data Input
                                                 .ENA(ena[12]),    // Port A RAM Enable Input
                                                 .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                 .WEA(wea),         // Port A Write Enable Input
                                                 .CLKB(clkb),      // Port B Clock
                                                 .DOB(doutb[102]),  // Port B 1-bit Data Output
                                                 .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                 .DIB(dinb[102]),   // Port B 1-bit Data Input
                                                 .ENB(enb[12]),    // Port B RAM Enable Input
                                                 .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                 .WEB(web)         // Port B Write Enable Input
                                                 ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_103 (
                                                 .CLKA(clka),      // Port A Clock
                                                 .DOA(douta[103]),  // Port A 1-bit Data Output
                                                 .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                 .DIA(dina[103]),   // Port A 1-bit Data Input
                                                 .ENA(ena[12]),    // Port A RAM Enable Input
                                                 .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                 .WEA(wea),         // Port A Write Enable Input
                                                 .CLKB(clkb),      // Port B Clock
                                                 .DOB(doutb[103]),  // Port B 1-bit Data Output
                                                 .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                 .DIB(dinb[103]),   // Port B 1-bit Data Input
                                                 .ENB(enb[12]),    // Port B RAM Enable Input
                                                 .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                 .WEB(web)         // Port B Write Enable Input
                                                 ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_104 (
                                                 .CLKA(clka),      // Port A Clock
                                                 .DOA(douta[104]),  // Port A 1-bit Data Output
                                                 .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                 .DIA(dina[104]),   // Port A 1-bit Data Input
                                                 .ENA(ena[13]),    // Port A RAM Enable Input
                                                 .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                 .WEA(wea),         // Port A Write Enable Input
                                                 .CLKB(clkb),      // Port B Clock
                                                 .DOB(doutb[104]),  // Port B 1-bit Data Output
                                                 .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                 .DIB(dinb[104]),   // Port B 1-bit Data Input
                                                 .ENB(enb[13]),    // Port B RAM Enable Input
                                                 .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                 .WEB(web)         // Port B Write Enable Input
                                                 ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_105 (
                                                 .CLKA(clka),      // Port A Clock
                                                 .DOA(douta[105]),  // Port A 1-bit Data Output
                                                 .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                 .DIA(dina[105]),   // Port A 1-bit Data Input
                                                 .ENA(ena[13]),    // Port A RAM Enable Input
                                                 .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                 .WEA(wea),         // Port A Write Enable Input
                                                 .CLKB(clkb),      // Port B Clock
                                                 .DOB(doutb[105]),  // Port B 1-bit Data Output
                                                 .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                 .DIB(dinb[105]),   // Port B 1-bit Data Input
                                                 .ENB(enb[13]),    // Port B RAM Enable Input
                                                 .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                 .WEB(web)         // Port B Write Enable Input
                                                 ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_106 (
                                                 .CLKA(clka),      // Port A Clock
                                                 .DOA(douta[106]),  // Port A 1-bit Data Output
                                                 .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                 .DIA(dina[106]),   // Port A 1-bit Data Input
                                                 .ENA(ena[13]),    // Port A RAM Enable Input
                                                 .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                 .WEA(wea),         // Port A Write Enable Input
                                                 .CLKB(clkb),      // Port B Clock
                                                 .DOB(doutb[106]),  // Port B 1-bit Data Output
                                                 .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                 .DIB(dinb[106]),   // Port B 1-bit Data Input
                                                 .ENB(enb[13]),    // Port B RAM Enable Input
                                                 .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                 .WEB(web)         // Port B Write Enable Input
                                                 ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_107 (
                                                 .CLKA(clka),      // Port A Clock
                                                 .DOA(douta[107]),  // Port A 1-bit Data Output
                                                 .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                 .DIA(dina[107]),   // Port A 1-bit Data Input
                                                 .ENA(ena[13]),    // Port A RAM Enable Input
                                                 .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                 .WEA(wea),         // Port A Write Enable Input
                                                 .CLKB(clkb),      // Port B Clock
                                                 .DOB(doutb[107]),  // Port B 1-bit Data Output
                                                 .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                 .DIB(dinb[107]),   // Port B 1-bit Data Input
                                                 .ENB(enb[13]),    // Port B RAM Enable Input
                                                 .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                 .WEB(web)         // Port B Write Enable Input
                                                 ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_108 (
                                                 .CLKA(clka),      // Port A Clock
                                                 .DOA(douta[108]),  // Port A 1-bit Data Output
                                                 .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                 .DIA(dina[108]),   // Port A 1-bit Data Input
                                                 .ENA(ena[13]),    // Port A RAM Enable Input
                                                 .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                 .WEA(wea),         // Port A Write Enable Input
                                                 .CLKB(clkb),      // Port B Clock
                                                 .DOB(doutb[108]),  // Port B 1-bit Data Output
                                                 .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                 .DIB(dinb[108]),   // Port B 1-bit Data Input
                                                 .ENB(enb[13]),    // Port B RAM Enable Input
                                                 .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                 .WEB(web)         // Port B Write Enable Input
                                                 ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_109 (
                                                 .CLKA(clka),      // Port A Clock
                                                 .DOA(douta[109]),  // Port A 1-bit Data Output
                                                 .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                 .DIA(dina[109]),   // Port A 1-bit Data Input
                                                 .ENA(ena[13]),    // Port A RAM Enable Input
                                                 .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                 .WEA(wea),         // Port A Write Enable Input
                                                 .CLKB(clkb),      // Port B Clock
                                                 .DOB(doutb[109]),  // Port B 1-bit Data Output
                                                 .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                 .DIB(dinb[109]),   // Port B 1-bit Data Input
                                                 .ENB(enb[13]),    // Port B RAM Enable Input
                                                 .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                 .WEB(web)         // Port B Write Enable Input
                                                 ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_110 (
                                                 .CLKA(clka),      // Port A Clock
                                                 .DOA(douta[110]),  // Port A 1-bit Data Output
                                                 .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                 .DIA(dina[110]),   // Port A 1-bit Data Input
                                                 .ENA(ena[13]),    // Port A RAM Enable Input
                                                 .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                 .WEA(wea),         // Port A Write Enable Input
                                                 .CLKB(clkb),      // Port B Clock
                                                 .DOB(doutb[110]),  // Port B 1-bit Data Output
                                                 .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                 .DIB(dinb[110]),   // Port B 1-bit Data Input
                                                 .ENB(enb[13]),    // Port B RAM Enable Input
                                                 .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                 .WEB(web)         // Port B Write Enable Input
                                                 ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_111 (
                                                 .CLKA(clka),      // Port A Clock
                                                 .DOA(douta[111]),  // Port A 1-bit Data Output
                                                 .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                 .DIA(dina[111]),   // Port A 1-bit Data Input
                                                 .ENA(ena[13]),    // Port A RAM Enable Input
                                                 .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                 .WEA(wea),         // Port A Write Enable Input
                                                 .CLKB(clkb),      // Port B Clock
                                                 .DOB(doutb[111]),  // Port B 1-bit Data Output
                                                 .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                 .DIB(dinb[111]),   // Port B 1-bit Data Input
                                                 .ENB(enb[13]),    // Port B RAM Enable Input
                                                 .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                 .WEB(web)         // Port B Write Enable Input
                                                 ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_112 (
                                                 .CLKA(clka),      // Port A Clock
                                                 .DOA(douta[112]),  // Port A 1-bit Data Output
                                                 .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                 .DIA(dina[112]),   // Port A 1-bit Data Input
                                                 .ENA(ena[14]),    // Port A RAM Enable Input
                                                 .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                 .WEA(wea),         // Port A Write Enable Input
                                                 .CLKB(clkb),      // Port B Clock
                                                 .DOB(doutb[112]),  // Port B 1-bit Data Output
                                                 .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                 .DIB(dinb[112]),   // Port B 1-bit Data Input
                                                 .ENB(enb[14]),    // Port B RAM Enable Input
                                                 .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                 .WEB(web)         // Port B Write Enable Input
                                                 ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_113 (
                                                 .CLKA(clka),      // Port A Clock
                                                 .DOA(douta[113]),  // Port A 1-bit Data Output
                                                 .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                 .DIA(dina[113]),   // Port A 1-bit Data Input
                                                 .ENA(ena[14]),    // Port A RAM Enable Input
                                                 .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                 .WEA(wea),         // Port A Write Enable Input
                                                 .CLKB(clkb),      // Port B Clock
                                                 .DOB(doutb[113]),  // Port B 1-bit Data Output
                                                 .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                 .DIB(dinb[113]),   // Port B 1-bit Data Input
                                                 .ENB(enb[14]),    // Port B RAM Enable Input
                                                 .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                 .WEB(web)         // Port B Write Enable Input
                                                 ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_114 (
                                                 .CLKA(clka),      // Port A Clock
                                                 .DOA(douta[114]),  // Port A 1-bit Data Output
                                                 .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                 .DIA(dina[114]),   // Port A 1-bit Data Input
                                                 .ENA(ena[14]),    // Port A RAM Enable Input
                                                 .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                 .WEA(wea),         // Port A Write Enable Input
                                                 .CLKB(clkb),      // Port B Clock
                                                 .DOB(doutb[114]),  // Port B 1-bit Data Output
                                                 .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                 .DIB(dinb[114]),   // Port B 1-bit Data Input
                                                 .ENB(enb[14]),    // Port B RAM Enable Input
                                                 .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                 .WEB(web)         // Port B Write Enable Input
                                                 ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_115 (
                                                 .CLKA(clka),      // Port A Clock
                                                 .DOA(douta[115]),  // Port A 1-bit Data Output
                                                 .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                 .DIA(dina[115]),   // Port A 1-bit Data Input
                                                 .ENA(ena[14]),    // Port A RAM Enable Input
                                                 .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                 .WEA(wea),         // Port A Write Enable Input
                                                 .CLKB(clkb),      // Port B Clock
                                                 .DOB(doutb[115]),  // Port B 1-bit Data Output
                                                 .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                 .DIB(dinb[115]),   // Port B 1-bit Data Input
                                                 .ENB(enb[14]),    // Port B RAM Enable Input
                                                 .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                 .WEB(web)         // Port B Write Enable Input
                                                 ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_116 (
                                                 .CLKA(clka),      // Port A Clock
                                                 .DOA(douta[116]),  // Port A 1-bit Data Output
                                                 .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                 .DIA(dina[116]),   // Port A 1-bit Data Input
                                                 .ENA(ena[14]),    // Port A RAM Enable Input
                                                 .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                 .WEA(wea),         // Port A Write Enable Input
                                                 .CLKB(clkb),      // Port B Clock
                                                 .DOB(doutb[116]),  // Port B 1-bit Data Output
                                                 .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                 .DIB(dinb[116]),   // Port B 1-bit Data Input
                                                 .ENB(enb[14]),    // Port B RAM Enable Input
                                                 .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                 .WEB(web)         // Port B Write Enable Input
                                                 ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_117 (
                                                 .CLKA(clka),      // Port A Clock
                                                 .DOA(douta[117]),  // Port A 1-bit Data Output
                                                 .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                 .DIA(dina[117]),   // Port A 1-bit Data Input
                                                 .ENA(ena[14]),    // Port A RAM Enable Input
                                                 .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                 .WEA(wea),         // Port A Write Enable Input
                                                 .CLKB(clkb),      // Port B Clock
                                                 .DOB(doutb[117]),  // Port B 1-bit Data Output
                                                 .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                 .DIB(dinb[117]),   // Port B 1-bit Data Input
                                                 .ENB(enb[14]),    // Port B RAM Enable Input
                                                 .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                 .WEB(web)         // Port B Write Enable Input
                                                 ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_118 (
                                                 .CLKA(clka),      // Port A Clock
                                                 .DOA(douta[118]),  // Port A 1-bit Data Output
                                                 .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                 .DIA(dina[118]),   // Port A 1-bit Data Input
                                                 .ENA(ena[14]),    // Port A RAM Enable Input
                                                 .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                 .WEA(wea),         // Port A Write Enable Input
                                                 .CLKB(clkb),      // Port B Clock
                                                 .DOB(doutb[118]),  // Port B 1-bit Data Output
                                                 .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                 .DIB(dinb[118]),   // Port B 1-bit Data Input
                                                 .ENB(enb[14]),    // Port B RAM Enable Input
                                                 .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                 .WEB(web)         // Port B Write Enable Input
                                                 ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_119 (
                                                 .CLKA(clka),      // Port A Clock
                                                 .DOA(douta[119]),  // Port A 1-bit Data Output
                                                 .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                 .DIA(dina[119]),   // Port A 1-bit Data Input
                                                 .ENA(ena[14]),    // Port A RAM Enable Input
                                                 .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                 .WEA(wea),         // Port A Write Enable Input
                                                 .CLKB(clkb),      // Port B Clock
                                                 .DOB(doutb[119]),  // Port B 1-bit Data Output
                                                 .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                 .DIB(dinb[119]),   // Port B 1-bit Data Input
                                                 .ENB(enb[14]),    // Port B RAM Enable Input
                                                 .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                 .WEB(web)         // Port B Write Enable Input
                                                 ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_120 (
                                                 .CLKA(clka),      // Port A Clock
                                                 .DOA(douta[120]),  // Port A 1-bit Data Output
                                                 .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                 .DIA(dina[120]),   // Port A 1-bit Data Input
                                                 .ENA(ena[15]),    // Port A RAM Enable Input
                                                 .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                 .WEA(wea),         // Port A Write Enable Input
                                                 .CLKB(clkb),      // Port B Clock
                                                 .DOB(doutb[120]),  // Port B 1-bit Data Output
                                                 .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                 .DIB(dinb[120]),   // Port B 1-bit Data Input
                                                 .ENB(enb[15]),    // Port B RAM Enable Input
                                                 .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                 .WEB(web)         // Port B Write Enable Input
                                                 ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_121 (
                                                 .CLKA(clka),      // Port A Clock
                                                 .DOA(douta[121]),  // Port A 1-bit Data Output
                                                 .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                 .DIA(dina[121]),   // Port A 1-bit Data Input
                                                 .ENA(ena[15]),    // Port A RAM Enable Input
                                                 .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                 .WEA(wea),         // Port A Write Enable Input
                                                 .CLKB(clkb),      // Port B Clock
                                                 .DOB(doutb[121]),  // Port B 1-bit Data Output
                                                 .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                 .DIB(dinb[121]),   // Port B 1-bit Data Input
                                                 .ENB(enb[15]),    // Port B RAM Enable Input
                                                 .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                 .WEB(web)         // Port B Write Enable Input
                                                 ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_122 (
                                                 .CLKA(clka),      // Port A Clock
                                                 .DOA(douta[122]),  // Port A 1-bit Data Output
                                                 .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                 .DIA(dina[122]),   // Port A 1-bit Data Input
                                                 .ENA(ena[15]),    // Port A RAM Enable Input
                                                 .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                 .WEA(wea),         // Port A Write Enable Input
                                                 .CLKB(clkb),      // Port B Clock
                                                 .DOB(doutb[122]),  // Port B 1-bit Data Output
                                                 .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                 .DIB(dinb[122]),   // Port B 1-bit Data Input
                                                 .ENB(enb[15]),    // Port B RAM Enable Input
                                                 .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                 .WEB(web)         // Port B Write Enable Input
                                                 ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_123 (
                                                 .CLKA(clka),      // Port A Clock
                                                 .DOA(douta[123]),  // Port A 1-bit Data Output
                                                 .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                 .DIA(dina[123]),   // Port A 1-bit Data Input
                                                 .ENA(ena[15]),    // Port A RAM Enable Input
                                                 .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                 .WEA(wea),         // Port A Write Enable Input
                                                 .CLKB(clkb),      // Port B Clock
                                                 .DOB(doutb[123]),  // Port B 1-bit Data Output
                                                 .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                 .DIB(dinb[123]),   // Port B 1-bit Data Input
                                                 .ENB(enb[15]),    // Port B RAM Enable Input
                                                 .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                 .WEB(web)         // Port B Write Enable Input
                                                 ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_124 (
                                                 .CLKA(clka),      // Port A Clock
                                                 .DOA(douta[124]),  // Port A 1-bit Data Output
                                                 .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                 .DIA(dina[124]),   // Port A 1-bit Data Input
                                                 .ENA(ena[15]),    // Port A RAM Enable Input
                                                 .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                 .WEA(wea),         // Port A Write Enable Input
                                                 .CLKB(clkb),      // Port B Clock
                                                 .DOB(doutb[124]),  // Port B 1-bit Data Output
                                                 .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                 .DIB(dinb[124]),   // Port B 1-bit Data Input
                                                 .ENB(enb[15]),    // Port B RAM Enable Input
                                                 .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                 .WEB(web)         // Port B Write Enable Input
                                                 ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_125 (
                                                 .CLKA(clka),      // Port A Clock
                                                 .DOA(douta[125]),  // Port A 1-bit Data Output
                                                 .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                 .DIA(dina[125]),   // Port A 1-bit Data Input
                                                 .ENA(ena[15]),    // Port A RAM Enable Input
                                                 .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                 .WEA(wea),         // Port A Write Enable Input
                                                 .CLKB(clkb),      // Port B Clock
                                                 .DOB(doutb[125]),  // Port B 1-bit Data Output
                                                 .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                 .DIB(dinb[125]),   // Port B 1-bit Data Input
                                                 .ENB(enb[15]),    // Port B RAM Enable Input
                                                 .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                 .WEB(web)         // Port B Write Enable Input
                                                 ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_126 (
                                                 .CLKA(clka),      // Port A Clock
                                                 .DOA(douta[126]),  // Port A 1-bit Data Output
                                                 .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                 .DIA(dina[126]),   // Port A 1-bit Data Input
                                                 .ENA(ena[15]),    // Port A RAM Enable Input
                                                 .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                 .WEA(wea),         // Port A Write Enable Input
                                                 .CLKB(clkb),      // Port B Clock
                                                 .DOB(doutb[126]),  // Port B 1-bit Data Output
                                                 .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                 .DIB(dinb[126]),   // Port B 1-bit Data Input
                                                 .ENB(enb[15]),    // Port B RAM Enable Input
                                                 .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                 .WEB(web)         // Port B Write Enable Input
                                                 ); // 

   RAMB16_S1_S1 #(
                  ) RAMB16_S1_S1_inst_128_0_127 (
                                                 .CLKA(clka),      // Port A Clock
                                                 .DOA(douta[127]),  // Port A 1-bit Data Output
                                                 .ADDRA(addra[13:0]),    // Port A 14-bit Address Input
                                                 .DIA(dina[127]),   // Port A 1-bit Data Input
                                                 .ENA(ena[15]),    // Port A RAM Enable Input
                                                 .SSRA(1'b0),     // Port A Synchronous Set/Reset Input
                                                 .WEA(wea),         // Port A Write Enable Input
                                                 .CLKB(clkb),      // Port B Clock
                                                 .DOB(doutb[127]),  // Port B 1-bit Data Output
                                                 .ADDRB(addrb[13:0]),    // Port B 14-bit Address Input
                                                 .DIB(dinb[127]),   // Port B 1-bit Data Input
                                                 .ENB(enb[15]),    // Port B RAM Enable Input
                                                 .SSRB(1'b0),     // Port B Synchronous Set/Reset Input
                                                 .WEB(web)         // Port B Write Enable Input
                                                 ); // 

endmodule
